module Controller
(input clk,
input [5:0] Opcode, Funct,
output MemToReg, RegDst, IorD, PCSrc, ALUSrcA, ALUSrcB, IRWrite, MemWrite, PCWrite, Branch, RegWrite, ALUControl
);

//implement FSM here



endmodule